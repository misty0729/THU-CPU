        "0110100100000001", -- LI R1 1;
		"0110101000000001", -- LI R2 1;
		"0110101110000101", -- LI R3 85;
		"0011001101100000", -- SLL R3 R3 0;
		"0110110000000101", -- LI R4 5;
		"1101101100100000", -- SW R3 R1 0;
		"0100100100000010", -- ADDIU R1 2;
		"0100101100000001", -- ADDIU R3 1;
		"0100110011111111", -- ADDIU R4 FF;
		"0010110011111100", -- BNEZ R4 Fc